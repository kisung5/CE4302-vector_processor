// Vector load/store unit

module vector_ldst #(parameter N = 32, V = 128) (
);


endmodule 
// MOV module
module mov_vector #(V = 128, N = 32)
(
input logic [V-1:0] inm
);

endmodule 